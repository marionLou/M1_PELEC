
module qbert_test2 (
	button_external_connection_export,
	clk_clk,
	reset_reset_n,
	switches_external_connection_export);	

	input		button_external_connection_export;
	input		clk_clk;
	input		reset_reset_n;
	input	[3:0]	switches_external_connection_export;
endmodule
